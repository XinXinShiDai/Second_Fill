module Reduce(
input [7:0] Din,
output Dout
    );

assign Dout = Din[0];

endmodule